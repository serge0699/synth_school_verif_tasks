// TODO: create interface

    // interface inv_if(input logic clk);
    // ..
    // endinterface

// Interface must contain single-bit logic fields:
// signal_in and signal_out
