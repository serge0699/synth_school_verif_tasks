// TODO: create cfg class

    // class cfg;
    // ..
    // enclass

// Class must containt int fields:
// latency and amount with default values 1 and 100
