    class array_alu_checker_base;

        //

    endclass