// TODO: create transaction class

    // class transaction;
    // ..
    // enclass

// Class must containt single-bit bit fields:
// signal_in and signal_out
