module testbench;

    class base1;
        rand bit [7:0] a;
             bit [7:0] b;
    endclass 

    base1 b1;
    initial begin
        b1 = new();
        repeat(5) begin
            b1.randomize();
            $display("b1.a: %8b", b1.a);
            $display("b1.b: %8b", b1.b);
        end
    end

endmodule

