module testbench;


    // TODO:
    //
    // Создайте поля:
    //   - bit [7:0] a
    //   - bit [7:0] b
    //
    // Опишите ограничения такие, что:
    //   1) 'b' больше 0
    //   2) 'a' делится на 'b' без остатка
    //   3) 'a' больше 'b'
    //   4) сумма 'a' и 'b' больше 100

    class my_class_1;


    endclass


    // TODO:
    //
    // Создайте поля:
    //   - bit [7:0] a
    //   - bit [7:0] b
    //
    // Опишите ограничения такие, что:
    //   1) если 'a' равно нулю, то 'b' равно 100
    //   2) 'a' меньше 100
    //   3) 'b' больше 50


    class my_class_2;


    endclass


    // TODO:
    //
    // Создайте поля:
    //   - int data []
    //
    // Опишите ограничения такие, что:
    //   1) размер массива четный
    //   2) размер массива меньше 10
    //   3) каждый элемент массива меньше 200
    //   4) если индекс элемента четный - элемент тоже четный

    class my_class_3;


    endclass


    // TODO:
    //
    // Создайте поля:
    //   - bit [1:0] size;
    //   - bit [7:0] data [];
    //
    // Опишите ограничения такие, что:
    //   1) размер 'data' равен 'size'
    //   2) если 'size' равен 3, то все элементы 'data' равны 0,
    //      иначе каждый элемент 'data' уникален

    class my_class_4;


    endclass


    // TODO:
    //
    // Создайте поля:
    //   - bit [7:0] data;
    //   - bit [7:0] addr;
    //   - bit req;
    //   - bit we;
    //
    // Опишите ограничения такие, что:
    //   1) адрес выровнен по границе 4 байт (последние 2 бита равны 0)
    //   2) если 'req' равен 1, то 'data' в интервале от 100 до 200
    //   3) если 'req' и 'we' равны 1, то 'addr' меньше 128

    class my_class_5;


    endclass


    // TODO:
    //
    // Создайте поля:
    //   - bit [31:0] tdata  [];
    //   - bit        tid;
    //   - bit        tlast [];
    //
    // Опишите ограничения такие, что:
    //   1) размер 'tdata' равен размеру 'tlast'
    //   2) размеры 'tdata' и 'tlast' меньше 33
    //   3) размеры 'tdata' и 'tlast' кратны 8
    //   4) 'tlast', равный 1, появляется в массиве не
    //      чаще, чем раз в 4 значения

    class my_class_6;


    endclass

    `include "checker.svh"

endmodule
