package test_pkg;

    // Пакет

    `include "packet.sv"

    // Конфигурация тестового сценария

    `include "cfg.sv"

    // Покрытие
    
    `include "coverage.sv"

    // Генератор

    `include "gen.sv"

    // Драйвер

    `include "driver.sv"

    // Монитор

    `include "monitor.sv"

    // Агент

    `include "agent.sv"

    // Проверка

    `include "checker.sv"

    // Окружение

    `include "env.sv"

    // Тест

    `include "test.sv"
    
endpackage